//-- Constantes para definir los valores del divisor segun la
//-- frecuencia deseada


//-------------------- Frecuencias
//-- Megaherzios  MHz
`define F_4MHz 3
`define F_3MHz 4
`define F_2MHz 6
`define F_1MHz 12

//-- Kilohercios KHz
`define F_4KHz 3000
`define F_3KHz 4000
`define F_2KHz 6000
`define F_1KHz 12000

//-- Hertzios (Hz)
`define F_2Hz   6000000
`define F_1Hz   12000000


//------- Frecuencias para notas musicales
//-- Octava 0
`define DO    45977  //-- 261 Hz
`define RE    40816  //-- 294 Hz
`define MI    36364  //-- 330 Hz
`define FA    34384  //-- 349 Hz
`define SOL   30612  //-- 392 Hz
`define LA    27273  //-- 440 Hz
`define SI    24291  //-- 494 Hz

//-- Octava 1
`define DO_1  22989  //--  2 * 261 Hz



