//-----------------------------------------------------------------------------
//-- Constantes para el modulo de generacion de baudios para comunicaciones serie
//------------------------------------------------------------------------------
//-- (C) BQ. September 2015. Written by Juan Gonzalez (Obijuan)
//------------------------------------------------------------------------------

//-- Para la icestick el calculo es el siguiente:
//-- Divisor = 16000000 / BAUDIOS  (Y se redondea a numero entero)

//-- Valores de los divisores para conseguir estos BAUDIOS:

`define B115200 138
`define B57600  277
`define B38400  416

`define B19200  833
`define B9600   1666
`define B4800   3333
`define B2400   6666
`define B1200   13333
`define B600    26666
`define B300    53333





